wire [49:0] up_arrow [49:0];
assign up_arrow[0] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[1] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[2] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[3] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[4] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[5] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[6] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[7] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[8] = 50'b00000000000000000000000111100000000000000000000000;
assign up_arrow[9] = 50'b00000000000000000000001111110000000000000000000000;
assign up_arrow[10] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[11] = 50'b00000000000000000000111111111100000000000000000000;
assign up_arrow[12] = 50'b00000000000000000001111111111110000000000000000000;
assign up_arrow[13] = 50'b00000000000000000011111111111111000000000000000000;
assign up_arrow[14] = 50'b00000000000000000111111111111111100000000000000000;
assign up_arrow[15] = 50'b00000000000000001111111111111111110000000000000000;
assign up_arrow[16] = 50'b00000000000000011111111111111111111000000000000000;
assign up_arrow[17] = 50'b00000000000000111111111111111111111100000000000000;
assign up_arrow[18] = 50'b00000000000001111111111111111111111110000000000000;
assign up_arrow[19] = 50'b00000000000011111111111111111111111111000000000000;
assign up_arrow[20] = 50'b00000000000111111111011111111011111111100000000000;
assign up_arrow[21] = 50'b00000000001111111000011111111000011111110000000000;
assign up_arrow[22] = 50'b00000000011111110000011111111000001111111000000000;
assign up_arrow[23] = 50'b00000000111111100000011111111000000111111100000000;
assign up_arrow[24] = 50'b00000001111111000000011111111000000011111110000000;
assign up_arrow[25] = 50'b00000001111110000000011111111000000001111110000000;
assign up_arrow[26] = 50'b00000001111100000000011111111000000000111110000000;
assign up_arrow[27] = 50'b00000001111000000000011111111000000000011110000000;
assign up_arrow[28] = 50'b00000001110000000000011111111000000000001110000000;
assign up_arrow[29] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[30] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[31] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[32] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[33] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[34] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[35] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[36] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[37] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[38] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[39] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[40] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[41] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[42] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[43] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow[44] = 50'b00000000000000000000001111110000000000000000000000;
assign up_arrow[45] = 50'b00000000000000000000000111100000000000000000000000;
assign up_arrow[46] = 50'b00000000000000000000000011000000000000000000000000;
assign up_arrow[47] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[48] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow[49] = 50'b00000000000000000000000000000000000000000000000000;
wire [49:0] left_arrow [49:0];
assign left_arrow[0] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[1] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[2] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[3] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[4] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[5] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[6] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[7] = 50'b00000000000000000000000011111000000000000000000000;
assign left_arrow[8] = 50'b00000000000000000000000111111000000000000000000000;
assign left_arrow[9] = 50'b00000000000000000000001111111000000000000000000000;
assign left_arrow[10] = 50'b00000000000000000000011111110000000000000000000000;
assign left_arrow[11] = 50'b00000000000000000000111111100000000000000000000000;
assign left_arrow[12] = 50'b00000000000000000001111111000000000000000000000000;
assign left_arrow[13] = 50'b00000000000000000011111110000000000000000000000000;
assign left_arrow[14] = 50'b00000000000000000111111100000000000000000000000000;
assign left_arrow[15] = 50'b00000000000000001111111000000000000000000000000000;
assign left_arrow[16] = 50'b00000000000000011111110000000000000000000000000000;
assign left_arrow[17] = 50'b00000000000000111111100000000000000000000000000000;
assign left_arrow[18] = 50'b00000000000001111111100000000000000000000000000000;
assign left_arrow[19] = 50'b00000000000011111111100000000000000000000000000000;
assign left_arrow[20] = 50'b00000000000111111111000000000000000000000000000000;
assign left_arrow[21] = 50'b00000000001111111111111111111111111111111111000000;
assign left_arrow[22] = 50'b00000000011111111111111111111111111111111111100000;
assign left_arrow[23] = 50'b00000000111111111111111111111111111111111111110000;
assign left_arrow[24] = 50'b00000000111111111111111111111111111111111111111000;
assign left_arrow[25] = 50'b00000000111111111111111111111111111111111111111000;
assign left_arrow[26] = 50'b00000000111111111111111111111111111111111111110000;
assign left_arrow[27] = 50'b00000000011111111111111111111111111111111111100000;
assign left_arrow[28] = 50'b00000000001111111111111111111111111111111111000000;
assign left_arrow[29] = 50'b00000000000111111111000000000000000000000000000000;
assign left_arrow[30] = 50'b00000000000011111111100000000000000000000000000000;
assign left_arrow[31] = 50'b00000000000001111111100000000000000000000000000000;
assign left_arrow[32] = 50'b00000000000000111111100000000000000000000000000000;
assign left_arrow[33] = 50'b00000000000000011111110000000000000000000000000000;
assign left_arrow[34] = 50'b00000000000000001111111000000000000000000000000000;
assign left_arrow[35] = 50'b00000000000000000111111100000000000000000000000000;
assign left_arrow[36] = 50'b00000000000000000011111110000000000000000000000000;
assign left_arrow[37] = 50'b00000000000000000001111111000000000000000000000000;
assign left_arrow[38] = 50'b00000000000000000000111111100000000000000000000000;
assign left_arrow[39] = 50'b00000000000000000000011111110000000000000000000000;
assign left_arrow[40] = 50'b00000000000000000000001111111000000000000000000000;
assign left_arrow[41] = 50'b00000000000000000000000111111000000000000000000000;
assign left_arrow[42] = 50'b00000000000000000000000011111000000000000000000000;
assign left_arrow[43] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[44] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[45] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[46] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[47] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[48] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow[49] = 50'b00000000000000000000000000000000000000000000000000;
wire [49:0] right_arrow [49:0];
assign right_arrow[0] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[1] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[2] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[3] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[4] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[5] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[6] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[7] = 50'b00000000000000000000011111000000000000000000000000;
assign right_arrow[8] = 50'b00000000000000000000011111100000000000000000000000;
assign right_arrow[9] = 50'b00000000000000000000011111110000000000000000000000;
assign right_arrow[10] = 50'b00000000000000000000001111111000000000000000000000;
assign right_arrow[11] = 50'b00000000000000000000000111111100000000000000000000;
assign right_arrow[12] = 50'b00000000000000000000000011111110000000000000000000;
assign right_arrow[13] = 50'b00000000000000000000000001111111000000000000000000;
assign right_arrow[14] = 50'b00000000000000000000000000111111100000000000000000;
assign right_arrow[15] = 50'b00000000000000000000000000011111110000000000000000;
assign right_arrow[16] = 50'b00000000000000000000000000001111111000000000000000;
assign right_arrow[17] = 50'b00000000000000000000000000000111111100000000000000;
assign right_arrow[18] = 50'b00000000000000000000000000000111111110000000000000;
assign right_arrow[19] = 50'b00000000000000000000000000000111111111000000000000;
assign right_arrow[20] = 50'b00000000000000000000000000000011111111100000000000;
assign right_arrow[21] = 50'b00000011111111111111111111111111111111110000000000;
assign right_arrow[22] = 50'b00000111111111111111111111111111111111111000000000;
assign right_arrow[23] = 50'b00001111111111111111111111111111111111111100000000;
assign right_arrow[24] = 50'b00011111111111111111111111111111111111111100000000;
assign right_arrow[25] = 50'b00011111111111111111111111111111111111111100000000;
assign right_arrow[26] = 50'b00001111111111111111111111111111111111111100000000;
assign right_arrow[27] = 50'b00000111111111111111111111111111111111111000000000;
assign right_arrow[28] = 50'b00000011111111111111111111111111111111110000000000;
assign right_arrow[29] = 50'b00000000000000000000000000000011111111100000000000;
assign right_arrow[30] = 50'b00000000000000000000000000000111111111000000000000;
assign right_arrow[31] = 50'b00000000000000000000000000000111111110000000000000;
assign right_arrow[32] = 50'b00000000000000000000000000000111111100000000000000;
assign right_arrow[33] = 50'b00000000000000000000000000001111111000000000000000;
assign right_arrow[34] = 50'b00000000000000000000000000011111110000000000000000;
assign right_arrow[35] = 50'b00000000000000000000000000111111100000000000000000;
assign right_arrow[36] = 50'b00000000000000000000000001111111000000000000000000;
assign right_arrow[37] = 50'b00000000000000000000000011111110000000000000000000;
assign right_arrow[38] = 50'b00000000000000000000000111111100000000000000000000;
assign right_arrow[39] = 50'b00000000000000000000001111111000000000000000000000;
assign right_arrow[40] = 50'b00000000000000000000011111110000000000000000000000;
assign right_arrow[41] = 50'b00000000000000000000011111100000000000000000000000;
assign right_arrow[42] = 50'b00000000000000000000011111000000000000000000000000;
assign right_arrow[43] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[44] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[45] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[46] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[47] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[48] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow[49] = 50'b00000000000000000000000000000000000000000000000000;
wire [49:0] down_arrow [49:0];
assign down_arrow[0] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[1] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[2] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[3] = 50'b00000000000000000000000011000000000000000000000000;
assign down_arrow[4] = 50'b00000000000000000000000111100000000000000000000000;
assign down_arrow[5] = 50'b00000000000000000000001111110000000000000000000000;
assign down_arrow[6] = 50'b00000000000000000000011111111000000000000000000000;
assign down_arrow[7] = 50'b00000000000000000000011111111100000000000000000000;
assign down_arrow[8] = 50'b00000000000000000000011111111100000000000000000000;
assign down_arrow[9] = 50'b00000000000000000000011111111100000000000000000000;
assign down_arrow[10] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[11] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[12] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[13] = 50'b0000000000000000000011111111100000000000000000000;
assign down_arrow[14] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[15] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[16] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[17] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[18] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[19] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[20] = 50'b00000000000000000000111111111000000000000000000000;
assign down_arrow[21] = 50'b00000001110000000000111111111000000000001110000000;
assign down_arrow[22] = 50'b00000001111000000000111111111000000000011110000000;
assign down_arrow[23] = 50'b00000001111100000000111111111000000000111110000000;
assign down_arrow[24] = 50'b00000001111110000000111111111000000001111110000000;
assign down_arrow[25] = 50'b00000001111111000000111111111000000011111110000000;
assign down_arrow[26] = 50'b00000000111111100000111111111000000111111100000000;
assign down_arrow[27] = 50'b00000000011111110000111111111000001111111000000000;
assign down_arrow[28] = 50'b00000000001111111000111111111000011111110000000000;
assign down_arrow[29] = 50'b00000000000111111111111111111011111111100000000000;
assign down_arrow[30] = 50'b00000000000011111111111111111111111111000000000000;
assign down_arrow[31] = 50'b00000000000001111111111111111111111110000000000000;
assign down_arrow[32] = 50'b00000000000000111111111111111111111100000000000000;
assign down_arrow[33] = 50'b00000000000000011111111111111111111000000000000000;
assign down_arrow[34] = 50'b00000000000000001111111111111111110000000000000000;
assign down_arrow[35] = 50'b00000000000000000111111111111111100000000000000000;
assign down_arrow[36] = 50'b00000000000000000011111111111111000000000000000000;
assign down_arrow[37] = 50'b00000000000000000001111111111110000000000000000000;
assign down_arrow[38] = 50'b00000000000000000000111111111100000000000000000000;
assign down_arrow[39] = 50'b00000000000000000000011111111000000000000000000000;
assign down_arrow[40] = 50'b00000000000000000000001111110000000000000000000000;
assign down_arrow[41] = 50'b00000000000000000000000111100000000000000000000000;
assign down_arrow[42] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[43] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[44] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[45] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[46] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[47] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[48] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow[49] = 50'b00000000000000000000000000000000000000000000000000;

wire [49:0] up_arrow_hollow [49:0];
assign up_arrow_hollow[0] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow_hollow[1] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow_hollow[2] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow_hollow[3] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow_hollow[4] = 50'b00000000000000000000000011000000000000000000000000;
assign up_arrow_hollow[5] = 50'b00000000000000000000000111100000000000000000000000;
assign up_arrow_hollow[6] = 50'b00000000000000000000001111110000000000000000000000;
assign up_arrow_hollow[7] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow_hollow[8] = 50'b00000000000000000000111100111100000000000000000000;
assign up_arrow_hollow[9] = 50'b00000000000000000001111000011110000000000000000000;
assign up_arrow_hollow[10] = 50'b00000000000000000011110000001111000000000000000000;
assign up_arrow_hollow[11] = 50'b00000000000000000111100000000111100000000000000000;
assign up_arrow_hollow[12] = 50'b00000000000000001111000000000011110000000000000000;
assign up_arrow_hollow[13] = 50'b00000000000000011110000000000001111000000000000000;
assign up_arrow_hollow[14] = 50'b00000000000000111100000000000000111100000000000000;
assign up_arrow_hollow[15] = 50'b00000000000001111000000000000000011110000000000000;
assign up_arrow_hollow[16] = 50'b00000000000011110000000010000000001111000000000000;
assign up_arrow_hollow[17] = 50'b00000000000111100000000111000000000111100000000000;
assign up_arrow_hollow[18] = 50'b00000000001111000000001111100000000011110000000000;
assign up_arrow_hollow[19] = 50'b00000000011110000000011000110000000001111000000000;
assign up_arrow_hollow[20] = 50'b00000000111100000011110000011111000000111100000000;
assign up_arrow_hollow[21] = 50'b00000001111000000111110000001111100000011110000000;
assign up_arrow_hollow[22] = 50'b00000011110000001111110000001111110000001111000000;
assign up_arrow_hollow[23] = 50'b00000111100000011111110000001111111000000111100000;
assign up_arrow_hollow[24] = 50'b00001111000000111111110000001111111100000011110000;
assign up_arrow_hollow[25] = 50'b00011110000001111011110000001110011110000011111000;
assign up_arrow_hollow[26] = 50'b00111110000011110011110000001110001111000011111000;
assign up_arrow_hollow[27] = 50'b00111110000111100011110000001110000111100011111100;
assign up_arrow_hollow[28] = 50'b00111111111111000011110011001110000011111111111000;
assign up_arrow_hollow[29] = 50'b00011111111110000011110111101110000001111111111000;
assign up_arrow_hollow[30] = 50'b00011111111100000001111000111110000000111111111000;
assign up_arrow_hollow[31] = 50'b00001111111000000001110000011110000000011111110000;
assign up_arrow_hollow[32] = 50'b00000111110000000001110000001110000000001111000000;
assign up_arrow_hollow[33] = 50'b00000000000000000011110000001110000000000000000000;
assign up_arrow_hollow[34] = 50'b00000000000000000011110000001110000000000000000000;
assign up_arrow_hollow[35] = 50'b00000000000000000011110000001110000000000000000000;
assign up_arrow_hollow[36] = 50'b00000000000000000011110000001110000000000000000000;
assign up_arrow_hollow[37] = 50'b00000000000000000011110000001110000000000000000000;
assign up_arrow_hollow[38] = 50'b00000000000000000011110000001110000000000000000000;
assign up_arrow_hollow[39] = 50'b00000000000000000011111000011110000000000000000000;
assign up_arrow_hollow[40] = 50'b00000000000000000011111100111110000000000000000000;
assign up_arrow_hollow[41] = 50'b00000000000000000001111111111110000000000000000000;
assign up_arrow_hollow[42] = 50'b00000000000000000000111111111100000000000000000000;
assign up_arrow_hollow[43] = 50'b00000000000000000000011111111000000000000000000000;
assign up_arrow_hollow[44] = 50'b00000000000000000000001111110000000000000000000000;
assign up_arrow_hollow[45] = 50'b00000000000000000000000111100000000000000000000000;
assign up_arrow_hollow[46] = 50'b00000000000000000000000011000000000000000000000000;
assign up_arrow_hollow[47] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow_hollow[48] = 50'b00000000000000000000000000000000000000000000000000;
assign up_arrow_hollow[49] = 50'b00000000000000000000000000000000000000000000000000;
wire [49:0] left_arrow_hollow [49:0];
assign left_arrow_hollow[0] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow_hollow[1] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow_hollow[2] = 50'b00000000000000000000000000010000000000000000000000;
assign left_arrow_hollow[3] = 50'b00000000000000000000000001111110000000000000000000;
assign left_arrow_hollow[4] = 50'b00000000000000000000000011111111000000000000000000;
assign left_arrow_hollow[5] = 50'b00000000000000000000000111111111000000000000000000;
assign left_arrow_hollow[6] = 50'b00000000000000000000001111111111100000000000000000;
assign left_arrow_hollow[7] = 50'b00000000000000000000011111111111100000000000000000;
assign left_arrow_hollow[8] = 50'b00000000000000000000111100001111100000000000000000;
assign left_arrow_hollow[9] = 50'b00000000000000000001111000001111100000000000000000;
assign left_arrow_hollow[10] = 50'b00000000000000000011110000001111000000000000000000;
assign left_arrow_hollow[11] = 50'b00000000000000000111100000011110000000000000000000;
assign left_arrow_hollow[12] = 50'b00000000000000001111000000111100000000000000000000;
assign left_arrow_hollow[13] = 50'b00000000000000011110000001111000000000000000000000;
assign left_arrow_hollow[14] = 50'b00000000000000111100000011110000000000000000000000;
assign left_arrow_hollow[15] = 50'b00000000000001111000000111100000000000000000000000;
assign left_arrow_hollow[16] = 50'b00000000000011110000001111000000000000000000000000;
assign left_arrow_hollow[17] = 50'b00000000000111100000011110000000000000000000000000;
assign left_arrow_hollow[18] = 50'b00000000001111000000111110000000000000000000000000;
assign left_arrow_hollow[19] = 50'b00000000011110000000111111111111111111111100000000;
assign left_arrow_hollow[20] = 50'b00000000111100000000111111111111111111111110000000;
assign left_arrow_hollow[21] = 50'b00000001111000000000111111111111111111111111000000;
assign left_arrow_hollow[22] = 50'b00000011110000000001100000000011000000011111100000;
assign left_arrow_hollow[23] = 50'b00000111100000000011000000000110000000001111110000;
assign left_arrow_hollow[24] = 50'b00001111000000000110000000001100000000000111111000;
assign left_arrow_hollow[25] = 50'b00001111000000001110000000001100000000000111111000;
assign left_arrow_hollow[26] = 50'b00000111100000000110000000000100000000001111110000;
assign left_arrow_hollow[27] = 50'b00000011110000000011000000000010000000011111100000;
assign left_arrow_hollow[28] = 50'b00000001111000000001111111111111111111111111000000;
assign left_arrow_hollow[29] = 50'b00000000111100000000111111111111111111111110000000;
assign left_arrow_hollow[30] = 50'b00000000011110000000111111111111111111111100000000;
assign left_arrow_hollow[31] = 50'b00000000001111000000111111111100011111111000000000;
assign left_arrow_hollow[32] = 50'b00000000000111100000011110000000000000000000000000;
assign left_arrow_hollow[33] = 50'b00000000000011110000001111000000000000000000000000;
assign left_arrow_hollow[34] = 50'b00000000000001111000000111100000000000000000000000;
assign left_arrow_hollow[35] = 50'b00000000000000111100000011110000000000000000000000;
assign left_arrow_hollow[36] = 50'b00000000000000011110000001111000000000000000000000;
assign left_arrow_hollow[37] = 50'b00000000000000001111000000111100000000000000000000;
assign left_arrow_hollow[38] = 50'b00000000000000000111100000011110000000000000000000;
assign left_arrow_hollow[39] = 50'b00000000000000000011110000001111000000000000000000;
assign left_arrow_hollow[40] = 50'b00000000000000000001111000001111100000000000000000;
assign left_arrow_hollow[41] = 50'b00000000000000000000111100001111100000000000000000;
assign left_arrow_hollow[42] = 50'b00000000000000000000011110001111100000000000000000;
assign left_arrow_hollow[43] = 50'b00000000000000000000001111111111100000000000000000;
assign left_arrow_hollow[44] = 50'b00000000000000000000000111111111100000000000000000;
assign left_arrow_hollow[45] = 50'b00000000000000000000000011111111000000000000000000;
assign left_arrow_hollow[46] = 50'b00000000000000000000000001111110000000000000000000;
assign left_arrow_hollow[47] = 50'b00000000000000000000000000111000000000000000000000;
assign left_arrow_hollow[48] = 50'b00000000000000000000000000000000000000000000000000;
assign left_arrow_hollow[49] = 50'b00000000000000000000000000000000000000000000000000;
wire [49:0] right_arrow_hollow [49:0];
assign right_arrow_hollow[0] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow_hollow[1] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow_hollow[2] = 50'b00000000000000000000011100000000000000000000000000;
assign right_arrow_hollow[3] = 50'b00000000000000000001111110000000000000000000000000;
assign right_arrow_hollow[4] = 50'b00000000000000000011111111000000000000000000000000;
assign right_arrow_hollow[5] = 50'b00000000000000000111111111100000000000000000000000;
assign right_arrow_hollow[6] = 50'b00000000000000000111111111110000000000000000000000;
assign right_arrow_hollow[7] = 50'b00000000000000000111110001111000000000000000000000;
assign right_arrow_hollow[8] = 50'b00000000000000000111110000111100000000000000000000;
assign right_arrow_hollow[9] = 50'b00000000000000000111110000011110000000000000000000;
assign right_arrow_hollow[10] = 50'b00000000000000000011110000001111000000000000000000;
assign right_arrow_hollow[11] = 50'b00000000000000000001111000000111100000000000000000;
assign right_arrow_hollow[12] = 50'b00000000000000000000111100000011110000000000000000;
assign right_arrow_hollow[13] = 50'b00000000000000000000011110000001111000000000000000;
assign right_arrow_hollow[14] = 50'b00000000000000000000001111000000111100000000000000;
assign right_arrow_hollow[15] = 50'b00000000000000000000000111100000011110000000000000;
assign right_arrow_hollow[16] = 50'b00000000000000000000000011110000001111000000000000;
assign right_arrow_hollow[17] = 50'b00000000000000000000000001111000000111100000000000;
assign right_arrow_hollow[18] = 50'b00000000011111111000111111111100000011110000000000;
assign right_arrow_hollow[19] = 50'b00000000111111111111111111111100000001111000000000;
assign right_arrow_hollow[20] = 50'b00000001111111111111111111111100000000111100000000;
assign right_arrow_hollow[21] = 50'b00000011111111111111111111111110000000011110000000;
assign right_arrow_hollow[22] = 50'b00000111111000000001000000000011000000001111000000;
assign right_arrow_hollow[23] = 50'b00001111110000000000100000000001100000000111100000;
assign right_arrow_hollow[24] = 50'b00011111100000000000110000000001110000000011110000;
assign right_arrow_hollow[25] = 50'b00011111100000000000110000000001100000000011110000;
assign right_arrow_hollow[26] = 50'b00001111110000000001100000000011000000000111100000;
assign right_arrow_hollow[27] = 50'b00000111111000000011000000000110000000001111000000;
assign right_arrow_hollow[28] = 50'b00000011111111111111111111111100000000011110000000;
assign right_arrow_hollow[29] = 50'b00000001111111111111111111111100000000111100000000;
assign right_arrow_hollow[30] = 50'b00000000111111111111111111111100000001111000000000;
assign right_arrow_hollow[31] = 50'b00000000000000000000000001111100000011110000000000;
assign right_arrow_hollow[32] = 50'b00000000000000000000000001111000000111100000000000;
assign right_arrow_hollow[33] = 50'b00000000000000000000000011110000001111000000000000;
assign right_arrow_hollow[34] = 50'b00000000000000000000000111100000011110000000000000;
assign right_arrow_hollow[35] = 50'b00000000000000000000001111000000111100000000000000;
assign right_arrow_hollow[36] = 50'b00000000000000000000011110000001111000000000000000;
assign right_arrow_hollow[37] = 50'b00000000000000000000111100000011110000000000000000;
assign right_arrow_hollow[38] = 50'b00000000000000000001111000000111100000000000000000;
assign right_arrow_hollow[39] = 50'b00000000000000000011110000001111000000000000000000;
assign right_arrow_hollow[40] = 50'b00000000000000000111110000011110000000000000000000;
assign right_arrow_hollow[41] = 50'b00000000000000000111110000111100000000000000000000;
assign right_arrow_hollow[42] = 50'b00000000000000000111111111111000000000000000000000;
assign right_arrow_hollow[43] = 50'b00000000000000000111111111110000000000000000000000;
assign right_arrow_hollow[44] = 50'b00000000000000000011111111100000000000000000000000;
assign right_arrow_hollow[45] = 50'b00000000000000000011111111000000000000000000000000;
assign right_arrow_hollow[46] = 50'b00000000000000000001111110000000000000000000000000;
assign right_arrow_hollow[47] = 50'b00000000000000000000001000000000000000000000000000;
assign right_arrow_hollow[48] = 50'b00000000000000000000000000000000000000000000000000;
assign right_arrow_hollow[49] = 50'b00000000000000000000000000000000000000000000000000;
wire [49:0] down_arrow_hollow [49:0];
assign down_arrow_hollow[0] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow_hollow[1] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow_hollow[2] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow_hollow[3] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow_hollow[4] = 50'b00000000000000000000000111100000000000000000000000;
assign down_arrow_hollow[5] = 50'b00000000000000000000001111110000000000000000000000;
assign down_arrow_hollow[6] = 50'b00000000000000000000011111111000000000000000000000;
assign down_arrow_hollow[7] = 50'b00000000000000000000111111111100000000000000000000;
assign down_arrow_hollow[8] = 50'b00000000000000000000111111111110000000000000000000;
assign down_arrow_hollow[9] = 50'b00000000000000000000111100111111000000000000000000;
assign down_arrow_hollow[10] = 50'b00000000000000000001111000011111000000000000000000;
assign down_arrow_hollow[11] = 50'b00000000000000000001110000001111000000000000000000;
assign down_arrow_hollow[12] = 50'b00000000000000000001110000001111000000000000000000;
assign down_arrow_hollow[13] = 50'b00000000000000000001110000001111000000000000000000;
assign down_arrow_hollow[14] = 50'b00000000000000000001110000001111000000000000000000;
assign down_arrow_hollow[15] = 50'b00000000000000000001110000001111000000000000000000;
assign down_arrow_hollow[16] = 50'b00000000000000000001110000001111000000000000000000;
assign down_arrow_hollow[17] = 50'b00000011110000000001110000001110000000001111100000;
assign down_arrow_hollow[18] = 50'b00001111111000000001111000001110000000011111110000;
assign down_arrow_hollow[19] = 50'b00011111111100000001111100011110000000111111111000;
assign down_arrow_hollow[20] = 50'b00011111111110000001110111101111000001111111111000;
assign down_arrow_hollow[21] = 50'b00011111111111000001110011001111000011111111111100;
assign down_arrow_hollow[22] = 50'b00111111000111100001110000001111000111100001111100;
assign down_arrow_hollow[23] = 50'b00011111000011110001110000001111001111000001111100;
assign down_arrow_hollow[24] = 50'b00011111000001111001110000001111011110000001111000;
assign down_arrow_hollow[25] = 50'b00001111000000111111110000001111111100000011110000;
assign down_arrow_hollow[26] = 50'b00000111100000011111110000001111111000000111100000;
assign down_arrow_hollow[27] = 50'b00000011110000001111110000001111110000001111000000;
assign down_arrow_hollow[28] = 50'b00000001111000000111110000001111100000011110000000;
assign down_arrow_hollow[29] = 50'b00000000111100000011111000001111000000111100000000;
assign down_arrow_hollow[30] = 50'b00000000011110000000001100011000000001111000000000;
assign down_arrow_hollow[31] = 50'b00000000001111000000000111110000000011110000000000;
assign down_arrow_hollow[32] = 50'b00000000000111100000000011100000000111100000000000;
assign down_arrow_hollow[33] = 50'b00000000000011110000000001000000001111000000000000;
assign down_arrow_hollow[34] = 50'b00000000000001111000000000000000011110000000000000;
assign down_arrow_hollow[35] = 50'b00000000000000111100000000000000111100000000000000;
assign down_arrow_hollow[36] = 50'b00000000000000011110000000000001111000000000000000;
assign down_arrow_hollow[37] = 50'b00000000000000001111000000000011110000000000000000;
assign down_arrow_hollow[38] = 50'b00000000000000000111100000000111100000000000000000;
assign down_arrow_hollow[39] = 50'b00000000000000000011110000001111000000000000000000;
assign down_arrow_hollow[40] = 50'b00000000000000000001111000011110000000000000000000;
assign down_arrow_hollow[41] = 50'b00000000000000000000111100111100000000000000000000;
assign down_arrow_hollow[42] = 50'b00000000000000000000011111111000000000000000000000;
assign down_arrow_hollow[43] = 50'b00000000000000000000001111110000000000000000000000;
assign down_arrow_hollow[44] = 50'b00000000000000000000000111100000000000000000000000;
assign down_arrow_hollow[45] = 50'b00000000000000000000000011000000000000000000000000;
assign down_arrow_hollow[46] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow_hollow[47] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow_hollow[48] = 50'b00000000000000000000000000000000000000000000000000;
assign down_arrow_hollow[49] = 50'b00000000000000000000000000000000000000000000000000;